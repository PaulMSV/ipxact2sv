
`define regmap0_addr_width 7
`define regmap0_data_width 8
